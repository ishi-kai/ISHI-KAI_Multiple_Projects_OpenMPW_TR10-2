* Created by KLayout

* cell OPAMP
* pin ib
* pin out
* pin vinn
* pin vdd
* pin vinp
* pin vss
.SUBCKT OPAMP 2 4 6 7 9 12
* net 2 ib
* net 4 out
* net 6 vinn
* net 7 vdd
* net 9 vinp
* net 12 vss
* device instance $1 r0 *1 -153.6,37.1 PMOS
M$1 7 2 1 7 PMOS L=5U W=30U AS=84P AD=45P PS=65.6U PD=33U
* device instance $2 r0 *1 -145.6,37.1 PMOS
M$2 2 2 7 7 PMOS L=5U W=30U AS=45P AD=84P PS=33U PD=65.6U
* device instance $3 r0 *1 -93.6,18.6 NMOS
M$3 10 10 12 12 NMOS L=5U W=120U AS=219P AD=180P PS=164.6U PD=132U
* device instance $7 r0 *1 -61.6,18.6 NMOS
M$7 5 10 12 12 NMOS L=5U W=120U AS=180P AD=219P PS=132U PD=164.6U
* device instance $11 m90 *1 151.3,122.6 PMOS
M$11 5 9 11 11 PMOS L=5U W=1080U AS=1698P AD=1698P PS=1196.6U PD=1196.6U
* device instance $29 r0 *1 -137.9,122.6 PMOS
M$29 10 6 11 11 PMOS L=5U W=1080U AS=1698P AD=1698P PS=1196.6U PD=1196.6U
* device instance $47 m0 *1 10.2,28.5 PMOS
M$47 4 2 7 7 PMOS L=5U W=600U AS=965P AD=965P PS=688.6U PD=688.6U
* device instance $59 m90 *1 127.3,38.3 NMOS
M$59 5 1 3 12 NMOS L=5U W=15U AS=42P AD=42P PS=35.6U PD=35.6U
* device instance $60 r90 *1 49.3,251 CSIO
C$60 4 3 12 8.856e-12 CSIO
* device instance $61 r270 *1 147,14.1 NMOS
M$61 4 5 12 12 NMOS L=5U W=200U AS=365P AD=365P PS=264.6U PD=264.6U
* device instance $65 r0 *1 -156.6,-4.8 NMOS
M$65 8 1 1 12 NMOS L=5U W=10U AS=28P AD=28P PS=25.6U PD=25.6U
* device instance $66 m90 *1 -143.6,-4.8 NMOS
M$66 8 8 12 12 NMOS L=5U W=10U AS=28P AD=28P PS=25.6U PD=25.6U
* device instance $67 r0 *1 -137.9,246.7 PMOS
M$67 11 2 7 7 PMOS L=5U W=720U AS=1158P AD=1158P PS=818.6U PD=818.6U
.ENDS OPAMP
