* Created by KLayout

* cell OPAMP_OHNO
* pin OUT
* pin VDD
* pin VSS
.SUBCKT OPAMP_OHNO 7 9 12
* net 7 OUT
* net 9 VDD
* net 12 VSS
* device instance $1 r0 *1 121.3,-48.2 NMOS
M$1 7 5 12 12 NMOS L=3U W=270U AS=444P AD=444P PS=329.6U PD=329.6U
* device instance $10 m135 *1 -63.8,-67.9 NMOS
M$10 5 3 2 12 NMOS L=3U W=30U AS=84P AD=84P PS=65.6U PD=65.6U
* device instance $11 m90 *1 -208.8,58.1 PMOS
M$11 3 1 9 9 PMOS L=3U W=120U AS=219P AD=219P PS=164.6U PD=164.6U
* device instance $15 r0 *1 -162.7,58.1 PMOS
M$15 6 1 9 9 PMOS L=3U W=240U AS=399P AD=399P PS=296.6U PD=296.6U
* device instance $23 r0 *1 -192.1,-59 NMOS
M$23 3 3 4 12 NMOS L=3U W=60U AS=129P AD=129P PS=98.6U PD=98.6U
* device instance $25 r0 *1 -227.7,-59 NMOS
M$25 4 4 12 12 NMOS L=3U W=60U AS=129P AD=129P PS=98.6U PD=98.6U
* device instance $27 r270 *1 -130.7,-29.8 NMOS
M$27 5 8 12 12 NMOS L=3U W=60U AS=129P AD=129P PS=98.6U PD=98.6U
* device instance $29 m45 *1 -130.7,-0.4 NMOS
M$29 8 8 12 12 NMOS L=3U W=60U AS=129P AD=129P PS=98.6U PD=98.6U
* device instance $31 m135 *1 -219.8,8.7 PMOS
M$31 1 1 9 9 PMOS L=3U W=90U AS=174P AD=174P PS=131.6U PD=131.6U
* device instance $34 m0 *1 121.3,14.1 PMOS
M$34 7 1 9 9 PMOS L=3U W=540U AS=888P AD=888P PS=659.2U PD=659.2U
* device instance $52 r0 *1 271.8,23.3 CSIO
C$52 7 2 12 8.856e-12 CSIO
* device instance $53 m0 *1 -74.5,-12.8 PMOS
M$53 5 10 6 6 PMOS L=3U W=720U AS=1158P AD=1158P PS=857.2U PD=857.2U
* device instance $77 r0 *1 -74.5,58.1 PMOS
M$77 8 11 6 6 PMOS L=3U W=720U AS=1158P AD=1158P PS=857.2U PD=857.2U
.ENDS OPAMP_OHNO
