** sch_path: /mnt/c/Data/OneDrive/MyDocuments/Community/ISHIKAI/shuttle/TR10/202509/OPAMP/opamp_matsushima/OPAMP_TR10-2-main/sch/opamp_cs_full.sch
.subckt opamp_cs_full vdd out vinp vinn vss
*.PININFO out:O vss:B vdd:B vinp:I vinn:I
XM1 vdd net1 net2 vdd PMOS w=13.6u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM2 net1 vinn net3 vss NMOS w=6.8u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM3 vdd net1 net1 vdd PMOS w=13.6u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM4 net2 vinp net3 vss NMOS w=6.8u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM5 vdd net5 net4 vdd PMOS w=27.2u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM6 vdd net5 net5 vdd PMOS w=27.2u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM7 net4 net4 vss vss NMOS w=20.4u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM8 net5 net5 vss vss NMOS w=20.4u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM9 net3 net4 vss vss NMOS w=3.4u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XM10 vdd net2 out vdd PMOS w=27.2u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
XC1 net2 out vss F_CSIO c=4p x=1u y=1u m=1
XM11 out net4 vss vss NMOS w=3.4u l=3.4u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 m=1
D2 vss vinp DN m=1
D1 vss vinn DN m=1
.ends
