* Created by KLayout

* cell OPAMP_matsushima
* pin out
* pin vdd
* pin vss
.SUBCKT OPAMP_matsushima 1 2 10
* net 1 out
* net 2 vdd
* net 10 vss
* device instance $1 r90 *1 23.1,-1.4 NDIO
D$1 10 8 NDIO A=12.96P P=14.4U
* device instance $2 r0 *1 -66.8,-1.1 NDIO
D$2 10 9 NDIO A=12.96P P=14.4U
* device instance $3 r270 *1 116.2,-6.3 CSIO
C$3 1 6 10 3.9952614e-12 CSIO
* device instance $4 m0 *1 -55.5,7.3 NMOS
M$4 7 9 5 10 NMOS L=3.4U W=6.8U AS=14.62P AD=14.62P PS=18.8U PD=18.8U
* device instance $6 r180 *1 11.8,7.1 NMOS
M$6 7 8 6 10 NMOS L=3.4U W=6.8U AS=14.62P AD=14.62P PS=18.8U PD=18.8U
* device instance $8 m0 *1 196.3,-51.3 NMOS
M$8 10 4 1 10 NMOS L=3.4U W=3.4U AS=9.52P AD=9.52P PS=12.4U PD=12.4U
* device instance $9 m0 *1 -4.9,-51.2 NMOS
M$9 10 4 7 10 NMOS L=3.4U W=3.4U AS=9.52P AD=9.52P PS=12.4U PD=12.4U
* device instance $10 r180 *1 -203.4,0.8 NMOS
M$10 10 3 3 10 NMOS L=3.4U W=20.4U AS=35.02P AD=35.02P PS=44.4U PD=44.4U
* device instance $16 r180 *1 -125.8,0.4 NMOS
M$16 10 4 4 10 NMOS L=3.4U W=20.4U AS=35.02P AD=35.02P PS=44.4U PD=44.4U
* device instance $22 m0 *1 190.5,54.1 PMOS
M$22 2 6 1 2 PMOS L=3.4U W=27.2U AS=45.22P AD=45.22P PS=57.2U PD=57.2U
* device instance $30 m0 *1 -168.8,39.4 PMOS
M$30 2 3 4 2 PMOS L=3.4U W=27.2U AS=45.22P AD=45.22P PS=57.2U PD=57.2U
* device instance $38 r180 *1 -206,39.4 PMOS
M$38 2 3 3 2 PMOS L=3.4U W=27.2U AS=45.22P AD=45.22P PS=57.2U PD=57.2U
* device instance $46 m0 *1 1.3,54.1 PMOS
M$46 2 5 6 2 PMOS L=3.4U W=13.6U AS=24.82P AD=24.82P PS=31.6U PD=31.6U
* device instance $50 r180 *1 -45.1,54.1 PMOS
M$50 2 5 5 2 PMOS L=3.4U W=13.6U AS=24.82P AD=24.82P PS=31.6U PD=31.6U
.ENDS OPAMP_matsushima
